module top_module(
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
);

    wire [15:0] w0, w1;
    wire sel;
    add16 inst1(.a(a[15:0]), .b(b[15:0]), .cin(1'b0), .cout(sel), .sum(sum[15:0]));
    add16 inst2(.a(a[31:16]), .b(b[31:16]), .cin(1'b0), .cout(), .sum(w0));
    add16 inst3(.a(a[31:16]), .b(b[31:16]), .cin(1'b1), .cout(), .sum(w1));
    
    assign sum[31:16] = sel ? w1:w0;
endmodule